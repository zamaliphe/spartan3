module systolic_PE6(inputword,outputword,clk30x, donext, reset);

`include "systolic_PE_core1.v"

`include "C_row6.v"

`include "systolic_PE_core2.v"

