module systolic_PE8(inputword,outputword,clk30x, donext, reset);

`include "systolic_PE_core1.v"

`include "C_row8.v"

`include "systolic_PE_core2.v"