module systolic_PE7(inputword,outputword,clk30x, donext, reset);

`include "systolic_PE_core1.v"

`include "C_row7.v"

`include "systolic_PE_core2.v"