module systolic_PE5(inputword,outputword,clk30x,donext, reset);

`include "systolic_PE_core1.v"

`include "C_row5.v"

`include "systolic_PE_core2.v"