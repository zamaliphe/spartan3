{begin template}
Ignore file {name}.vhd