library verilog;
use verilog.vl_types.all;
entity detailed_testbench is
end detailed_testbench;
