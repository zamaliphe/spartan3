library verilog;
use verilog.vl_types.all;
entity Transposer is
    generic(
        STEP_WIDTH      : integer := 3
    );
    port(
        transposer_clk  : in     vl_logic;
        transposer_reset: in     vl_logic;
        do_transpose    : in     vl_logic;
        do_bitreversing : in     vl_logic;
        done_transpose  : out    vl_logic;
        ram00_port0_add : out    vl_logic_vector(8 downto 0);
        ram00_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram00_port1_add : out    vl_logic_vector(8 downto 0);
        ram00_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram00_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram00_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram01_port0_add : out    vl_logic_vector(8 downto 0);
        ram01_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram01_port1_add : out    vl_logic_vector(8 downto 0);
        ram01_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram01_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram01_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram02_port0_add : out    vl_logic_vector(8 downto 0);
        ram02_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram02_port1_add : out    vl_logic_vector(8 downto 0);
        ram02_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram02_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram02_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram03_port0_add : out    vl_logic_vector(8 downto 0);
        ram03_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram03_port1_add : out    vl_logic_vector(8 downto 0);
        ram03_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram03_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram03_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram04_port0_add : out    vl_logic_vector(8 downto 0);
        ram04_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram04_port1_add : out    vl_logic_vector(8 downto 0);
        ram04_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram04_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram04_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram05_port0_add : out    vl_logic_vector(8 downto 0);
        ram05_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram05_port1_add : out    vl_logic_vector(8 downto 0);
        ram05_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram05_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram05_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram06_port0_add : out    vl_logic_vector(8 downto 0);
        ram06_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram06_port1_add : out    vl_logic_vector(8 downto 0);
        ram06_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram06_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram06_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram07_port0_add : out    vl_logic_vector(8 downto 0);
        ram07_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram07_port1_add : out    vl_logic_vector(8 downto 0);
        ram07_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram07_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram07_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram08_port0_add : out    vl_logic_vector(8 downto 0);
        ram08_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram08_port1_add : out    vl_logic_vector(8 downto 0);
        ram08_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram08_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram08_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram09_port0_add : out    vl_logic_vector(8 downto 0);
        ram09_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram09_port1_add : out    vl_logic_vector(8 downto 0);
        ram09_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram09_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram09_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram10_port0_add : out    vl_logic_vector(8 downto 0);
        ram10_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram10_port1_add : out    vl_logic_vector(8 downto 0);
        ram10_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram10_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram10_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram11_port0_add : out    vl_logic_vector(8 downto 0);
        ram11_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram11_port1_add : out    vl_logic_vector(8 downto 0);
        ram11_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram11_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram11_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram12_port0_add : out    vl_logic_vector(8 downto 0);
        ram12_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram12_port1_add : out    vl_logic_vector(8 downto 0);
        ram12_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram12_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram12_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram13_port0_add : out    vl_logic_vector(8 downto 0);
        ram13_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram13_port1_add : out    vl_logic_vector(8 downto 0);
        ram13_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram13_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram13_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram14_port0_add : out    vl_logic_vector(8 downto 0);
        ram14_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram14_port1_add : out    vl_logic_vector(8 downto 0);
        ram14_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram14_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram14_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram15_port0_add : out    vl_logic_vector(8 downto 0);
        ram15_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram15_port1_add : out    vl_logic_vector(8 downto 0);
        ram15_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram15_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram15_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram16_port0_add : out    vl_logic_vector(8 downto 0);
        ram16_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram16_port1_add : out    vl_logic_vector(8 downto 0);
        ram16_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram16_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram16_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram17_port0_add : out    vl_logic_vector(8 downto 0);
        ram17_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram17_port1_add : out    vl_logic_vector(8 downto 0);
        ram17_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram17_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram17_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram18_port0_add : out    vl_logic_vector(8 downto 0);
        ram18_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram18_port1_add : out    vl_logic_vector(8 downto 0);
        ram18_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram18_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram18_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram19_port0_add : out    vl_logic_vector(8 downto 0);
        ram19_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram19_port1_add : out    vl_logic_vector(8 downto 0);
        ram19_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram19_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram19_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram20_port0_add : out    vl_logic_vector(8 downto 0);
        ram20_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram20_port1_add : out    vl_logic_vector(8 downto 0);
        ram20_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram20_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram20_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram21_port0_add : out    vl_logic_vector(8 downto 0);
        ram21_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram21_port1_add : out    vl_logic_vector(8 downto 0);
        ram21_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram21_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram21_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram22_port0_add : out    vl_logic_vector(8 downto 0);
        ram22_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram22_port1_add : out    vl_logic_vector(8 downto 0);
        ram22_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram22_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram22_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram23_port0_add : out    vl_logic_vector(8 downto 0);
        ram23_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram23_port1_add : out    vl_logic_vector(8 downto 0);
        ram23_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram23_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram23_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram24_port0_add : out    vl_logic_vector(8 downto 0);
        ram24_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram24_port1_add : out    vl_logic_vector(8 downto 0);
        ram24_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram24_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram24_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram25_port0_add : out    vl_logic_vector(8 downto 0);
        ram25_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram25_port1_add : out    vl_logic_vector(8 downto 0);
        ram25_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram25_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram25_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram26_port0_add : out    vl_logic_vector(8 downto 0);
        ram26_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram26_port1_add : out    vl_logic_vector(8 downto 0);
        ram26_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram26_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram26_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram27_port0_add : out    vl_logic_vector(8 downto 0);
        ram27_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram27_port1_add : out    vl_logic_vector(8 downto 0);
        ram27_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram27_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram27_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram28_port0_add : out    vl_logic_vector(8 downto 0);
        ram28_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram28_port1_add : out    vl_logic_vector(8 downto 0);
        ram28_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram28_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram28_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram29_port0_add : out    vl_logic_vector(8 downto 0);
        ram29_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram29_port1_add : out    vl_logic_vector(8 downto 0);
        ram29_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram29_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram29_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram30_port0_add : out    vl_logic_vector(8 downto 0);
        ram30_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram30_port1_add : out    vl_logic_vector(8 downto 0);
        ram30_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram30_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram30_cs_we_oe_1: out    vl_logic_vector(2 downto 0);
        ram31_port0_add : out    vl_logic_vector(8 downto 0);
        ram31_port0_bus : inout  vl_logic_vector(15 downto 0);
        ram31_port1_add : out    vl_logic_vector(8 downto 0);
        ram31_port1_bus : inout  vl_logic_vector(15 downto 0);
        ram31_cs_we_oe_0: out    vl_logic_vector(2 downto 0);
        ram31_cs_we_oe_1: out    vl_logic_vector(2 downto 0)
    );
end Transposer;
