library verilog;
use verilog.vl_types.all;
entity detailed_testbench is
    generic(
        N               : integer := 4096
    );
end detailed_testbench;
