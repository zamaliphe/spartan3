library verilog;
use verilog.vl_types.all;
entity converter is
end converter;
