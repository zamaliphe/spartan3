library verilog;
use verilog.vl_types.all;
entity temp_MultTOP is
end temp_MultTOP;
