//Automatically generated using C code: Theja 2008
module Butterfly_Mult_Wallace(prod,a,b);
output[31:0] prod;
input[15:0] a,b;
wire p01;
wire p11;
wire p12;
wire p21;
wire p22;
wire p23;
wire p31;
wire p32;
wire p33;
wire p34;
wire p41;
wire p42;
wire p43;
wire p44;
wire p45;
wire p51;
wire p52;
wire p53;
wire p54;
wire p55;
wire p56;
wire p61;
wire p62;
wire p63;
wire p64;
wire p65;
wire p66;
wire p67;
wire p71;
wire p72;
wire p73;
wire p74;
wire p75;
wire p76;
wire p77;
wire p78;
wire p81;
wire p82;
wire p83;
wire p84;
wire p85;
wire p86;
wire p87;
wire p88;
wire p89;
wire p91;
wire p92;
wire p93;
wire p94;
wire p95;
wire p96;
wire p97;
wire p98;
wire p99;
wire p910;
wire p101;
wire p102;
wire p103;
wire p104;
wire p105;
wire p106;
wire p107;
wire p108;
wire p109;
wire p1010;
wire p1011;
wire p111;
wire p112;
wire p113;
wire p114;
wire p115;
wire p116;
wire p117;
wire p118;
wire p119;
wire p1110;
wire p1111;
wire p1112;
wire p121;
wire p122;
wire p123;
wire p124;
wire p125;
wire p126;
wire p127;
wire p128;
wire p129;
wire p1210;
wire p1211;
wire p1212;
wire p1213;
wire p131;
wire p132;
wire p133;
wire p134;
wire p135;
wire p136;
wire p137;
wire p138;
wire p139;
wire p1310;
wire p1311;
wire p1312;
wire p1313;
wire p1314;
wire p141;
wire p142;
wire p143;
wire p144;
wire p145;
wire p146;
wire p147;
wire p148;
wire p149;
wire p1410;
wire p1411;
wire p1412;
wire p1413;
wire p1414;
wire p1415;
wire p151;
wire p152;
wire p153;
wire p154;
wire p155;
wire p156;
wire p157;
wire p158;
wire p159;
wire p1510;
wire p1511;
wire p1512;
wire p1513;
wire p1514;
wire p1515;
wire p1516;
wire p301;
wire p291;
wire p292;
wire p281;
wire p282;
wire p283;
wire p271;
wire p272;
wire p273;
wire p274;
wire p261;
wire p262;
wire p263;
wire p264;
wire p265;
wire p251;
wire p252;
wire p253;
wire p254;
wire p255;
wire p256;
wire p241;
wire p242;
wire p243;
wire p244;
wire p245;
wire p246;
wire p247;
wire p231;
wire p232;
wire p233;
wire p234;
wire p235;
wire p236;
wire p237;
wire p238;
wire p221;
wire p222;
wire p223;
wire p224;
wire p225;
wire p226;
wire p227;
wire p228;
wire p229;
wire p211;
wire p212;
wire p213;
wire p214;
wire p215;
wire p216;
wire p217;
wire p218;
wire p219;
wire p2110;
wire p201;
wire p202;
wire p203;
wire p204;
wire p205;
wire p206;
wire p207;
wire p208;
wire p209;
wire p2010;
wire p2011;
wire p191;
wire p192;
wire p193;
wire p194;
wire p195;
wire p196;
wire p197;
wire p198;
wire p199;
wire p1910;
wire p1911;
wire p1912;
wire p181;
wire p182;
wire p183;
wire p184;
wire p185;
wire p186;
wire p187;
wire p188;
wire p189;
wire p1810;
wire p1811;
wire p1812;
wire p1813;
wire p171;
wire p172;
wire p173;
wire p174;
wire p175;
wire p176;
wire p177;
wire p178;
wire p179;
wire p1710;
wire p1711;
wire p1712;
wire p1713;
wire p1714;
wire p161;
wire p162;
wire p163;
wire p164;
wire p165;
wire p166;
wire p167;
wire p168;
wire p169;
wire p1610;
wire p1611;
wire p1612;
wire p1613;
wire p1614;
wire p1615;
wire[29:0] x;
wire[29:0] y;
wire[29:0] z;
wire t;
wire s1q17;
wire c1q17;
wire s1q16;
wire c1q16;
wire s1q15;
wire c1q15;
wire s1q14;
wire c1q14;
wire s2q18;
wire c2q18;
wire s2q17;
wire c2q17;
wire s2q16;
wire c2q16;
wire s2q15;
wire c2q15;
wire s2q14;
wire c2q14;
wire s2q13;
wire c2q13;
wire s3q19;
wire c3q19;
wire s3q18;
wire c3q18;
wire s3q17;
wire c3q17;
wire s3q16;
wire c3q16;
wire s3q15;
wire c3q15;
wire s3q14;
wire c3q14;
wire s3q13;
wire c3q13;
wire s3q12;
wire c3q12;
wire s4q20;
wire c4q20;
wire s4q19;
wire c4q19;
wire s4q18;
wire c4q18;
wire s4q17;
wire c4q17;
wire s4q16;
wire c4q16;
wire s4q15;
wire c4q15;
wire s4q14;
wire c4q14;
wire s4q13;
wire c4q13;
wire s4q12;
wire c4q12;
wire s4q11;
wire c4q11;
wire s5q21;
wire c5q21;
wire s5q20;
wire c5q20;
wire s5q19;
wire c5q19;
wire s5q18;
wire c5q18;
wire s5q17;
wire c5q17;
wire s5q16;
wire c5q16;
wire s5q15;
wire c5q15;
wire s5q14;
wire c5q14;
wire s5q13;
wire c5q13;
wire s5q12;
wire c5q12;
wire s5q11;
wire c5q11;
wire s5q10;
wire c5q10;
wire s6q22;
wire c6q22;
wire s6q21;
wire c6q21;
wire s6q20;
wire c6q20;
wire s6q19;
wire c6q19;
wire s6q18;
wire c6q18;
wire s6q17;
wire c6q17;
wire s6q16;
wire c6q16;
wire s6q15;
wire c6q15;
wire s6q14;
wire c6q14;
wire s6q13;
wire c6q13;
wire s6q12;
wire c6q12;
wire s6q11;
wire c6q11;
wire s6q10;
wire c6q10;
wire s6q9;
wire c6q9;
wire s7q23;
wire c7q23;
wire s7q22;
wire c7q22;
wire s7q21;
wire c7q21;
wire s7q20;
wire c7q20;
wire s7q19;
wire c7q19;
wire s7q18;
wire c7q18;
wire s7q17;
wire c7q17;
wire s7q16;
wire c7q16;
wire s7q15;
wire c7q15;
wire s7q14;
wire c7q14;
wire s7q13;
wire c7q13;
wire s7q12;
wire c7q12;
wire s7q11;
wire c7q11;
wire s7q10;
wire c7q10;
wire s7q9;
wire c7q9;
wire s7q8;
wire c7q8;
wire s8q24;
wire c8q24;
wire s8q23;
wire c8q23;
wire s8q22;
wire c8q22;
wire s8q21;
wire c8q21;
wire s8q20;
wire c8q20;
wire s8q19;
wire c8q19;
wire s8q18;
wire c8q18;
wire s8q17;
wire c8q17;
wire s8q16;
wire c8q16;
wire s8q15;
wire c8q15;
wire s8q14;
wire c8q14;
wire s8q13;
wire c8q13;
wire s8q12;
wire c8q12;
wire s8q11;
wire c8q11;
wire s8q10;
wire c8q10;
wire s8q9;
wire c8q9;
wire s8q8;
wire c8q8;
wire s8q7;
wire c8q7;
wire s9q25;
wire c9q25;
wire s9q24;
wire c9q24;
wire s9q23;
wire c9q23;
wire s9q22;
wire c9q22;
wire s9q21;
wire c9q21;
wire s9q20;
wire c9q20;
wire s9q19;
wire c9q19;
wire s9q18;
wire c9q18;
wire s9q17;
wire c9q17;
wire s9q16;
wire c9q16;
wire s9q15;
wire c9q15;
wire s9q14;
wire c9q14;
wire s9q13;
wire c9q13;
wire s9q12;
wire c9q12;
wire s9q11;
wire c9q11;
wire s9q10;
wire c9q10;
wire s9q9;
wire c9q9;
wire s9q8;
wire c9q8;
wire s9q7;
wire c9q7;
wire s9q6;
wire c9q6;
wire s10q26;
wire c10q26;
wire s10q25;
wire c10q25;
wire s10q24;
wire c10q24;
wire s10q23;
wire c10q23;
wire s10q22;
wire c10q22;
wire s10q21;
wire c10q21;
wire s10q20;
wire c10q20;
wire s10q19;
wire c10q19;
wire s10q18;
wire c10q18;
wire s10q17;
wire c10q17;
wire s10q16;
wire c10q16;
wire s10q15;
wire c10q15;
wire s10q14;
wire c10q14;
wire s10q13;
wire c10q13;
wire s10q12;
wire c10q12;
wire s10q11;
wire c10q11;
wire s10q10;
wire c10q10;
wire s10q9;
wire c10q9;
wire s10q8;
wire c10q8;
wire s10q7;
wire c10q7;
wire s10q6;
wire c10q6;
wire s10q5;
wire c10q5;
wire s11q27;
wire c11q27;
wire s11q26;
wire c11q26;
wire s11q25;
wire c11q25;
wire s11q24;
wire c11q24;
wire s11q23;
wire c11q23;
wire s11q22;
wire c11q22;
wire s11q21;
wire c11q21;
wire s11q20;
wire c11q20;
wire s11q19;
wire c11q19;
wire s11q18;
wire c11q18;
wire s11q17;
wire c11q17;
wire s11q16;
wire c11q16;
wire s11q15;
wire c11q15;
wire s11q14;
wire c11q14;
wire s11q13;
wire c11q13;
wire s11q12;
wire c11q12;
wire s11q11;
wire c11q11;
wire s11q10;
wire c11q10;
wire s11q9;
wire c11q9;
wire s11q8;
wire c11q8;
wire s11q7;
wire c11q7;
wire s11q6;
wire c11q6;
wire s11q5;
wire c11q5;
wire s11q4;
wire c11q4;
wire s12q28;
wire c12q28;
wire s12q27;
wire c12q27;
wire s12q26;
wire c12q26;
wire s12q25;
wire c12q25;
wire s12q24;
wire c12q24;
wire s12q23;
wire c12q23;
wire s12q22;
wire c12q22;
wire s12q21;
wire c12q21;
wire s12q20;
wire c12q20;
wire s12q19;
wire c12q19;
wire s12q18;
wire c12q18;
wire s12q17;
wire c12q17;
wire s12q16;
wire c12q16;
wire s12q15;
wire c12q15;
wire s12q14;
wire c12q14;
wire s12q13;
wire c12q13;
wire s12q12;
wire c12q12;
wire s12q11;
wire c12q11;
wire s12q10;
wire c12q10;
wire s12q9;
wire c12q9;
wire s12q8;
wire c12q8;
wire s12q7;
wire c12q7;
wire s12q6;
wire c12q6;
wire s12q5;
wire c12q5;
wire s12q4;
wire c12q4;
wire s12q3;
wire c12q3;
wire s13q29;
wire c13q29;
wire s13q28;
wire c13q28;
wire s13q27;
wire c13q27;
wire s13q26;
wire c13q26;
wire s13q25;
wire c13q25;
wire s13q24;
wire c13q24;
wire s13q23;
wire c13q23;
wire s13q22;
wire c13q22;
wire s13q21;
wire c13q21;
wire s13q20;
wire c13q20;
wire s13q19;
wire c13q19;
wire s13q18;
wire c13q18;
wire s13q17;
wire c13q17;
wire s13q16;
wire c13q16;
wire s13q15;
wire c13q15;
wire s13q14;
wire c13q14;
wire s13q13;
wire c13q13;
wire s13q12;
wire c13q12;
wire s13q11;
wire c13q11;
wire s13q10;
wire c13q10;
wire s13q9;
wire c13q9;
wire s13q8;
wire c13q8;
wire s13q7;
wire c13q7;
wire s13q6;
wire c13q6;
wire s13q5;
wire c13q5;
wire s13q4;
wire c13q4;
wire s13q3;
wire c13q3;
wire s13q2;
wire c13q2;
wire s1,s2,c1,c2;
and(p01,a[0],b[0]);
and(p11,a[1],b[0]);
and(p12,a[0],b[1]);
and(p21,a[2],b[0]);
and(p22,a[1],b[1]);
and(p23,a[0],b[2]);
and(p31,a[3],b[0]);
and(p32,a[2],b[1]);
and(p33,a[1],b[2]);
and(p34,a[0],b[3]);
and(p41,a[4],b[0]);
and(p42,a[3],b[1]);
and(p43,a[2],b[2]);
and(p44,a[1],b[3]);
and(p45,a[0],b[4]);
and(p51,a[5],b[0]);
and(p52,a[4],b[1]);
and(p53,a[3],b[2]);
and(p54,a[2],b[3]);
and(p55,a[1],b[4]);
and(p56,a[0],b[5]);
and(p61,a[6],b[0]);
and(p62,a[5],b[1]);
and(p63,a[4],b[2]);
and(p64,a[3],b[3]);
and(p65,a[2],b[4]);
and(p66,a[1],b[5]);
and(p67,a[0],b[6]);
and(p71,a[7],b[0]);
and(p72,a[6],b[1]);
and(p73,a[5],b[2]);
and(p74,a[4],b[3]);
and(p75,a[3],b[4]);
and(p76,a[2],b[5]);
and(p77,a[1],b[6]);
and(p78,a[0],b[7]);
and(p81,a[8],b[0]);
and(p82,a[7],b[1]);
and(p83,a[6],b[2]);
and(p84,a[5],b[3]);
and(p85,a[4],b[4]);
and(p86,a[3],b[5]);
and(p87,a[2],b[6]);
and(p88,a[1],b[7]);
and(p89,a[0],b[8]);
and(p91,a[9],b[0]);
and(p92,a[8],b[1]);
and(p93,a[7],b[2]);
and(p94,a[6],b[3]);
and(p95,a[5],b[4]);
and(p96,a[4],b[5]);
and(p97,a[3],b[6]);
and(p98,a[2],b[7]);
and(p99,a[1],b[8]);
and(p910,a[0],b[9]);
and(p101,a[10],b[0]);
and(p102,a[9],b[1]);
and(p103,a[8],b[2]);
and(p104,a[7],b[3]);
and(p105,a[6],b[4]);
and(p106,a[5],b[5]);
and(p107,a[4],b[6]);
and(p108,a[3],b[7]);
and(p109,a[2],b[8]);
and(p1010,a[1],b[9]);
and(p1011,a[0],b[10]);
and(p111,a[11],b[0]);
and(p112,a[10],b[1]);
and(p113,a[9],b[2]);
and(p114,a[8],b[3]);
and(p115,a[7],b[4]);
and(p116,a[6],b[5]);
and(p117,a[5],b[6]);
and(p118,a[4],b[7]);
and(p119,a[3],b[8]);
and(p1110,a[2],b[9]);
and(p1111,a[1],b[10]);
and(p1112,a[0],b[11]);
and(p121,a[12],b[0]);
and(p122,a[11],b[1]);
and(p123,a[10],b[2]);
and(p124,a[9],b[3]);
and(p125,a[8],b[4]);
and(p126,a[7],b[5]);
and(p127,a[6],b[6]);
and(p128,a[5],b[7]);
and(p129,a[4],b[8]);
and(p1210,a[3],b[9]);
and(p1211,a[2],b[10]);
and(p1212,a[1],b[11]);
and(p1213,a[0],b[12]);
and(p131,a[13],b[0]);
and(p132,a[12],b[1]);
and(p133,a[11],b[2]);
and(p134,a[10],b[3]);
and(p135,a[9],b[4]);
and(p136,a[8],b[5]);
and(p137,a[7],b[6]);
and(p138,a[6],b[7]);
and(p139,a[5],b[8]);
and(p1310,a[4],b[9]);
and(p1311,a[3],b[10]);
and(p1312,a[2],b[11]);
and(p1313,a[1],b[12]);
and(p1314,a[0],b[13]);
and(p141,a[14],b[0]);
and(p142,a[13],b[1]);
and(p143,a[12],b[2]);
and(p144,a[11],b[3]);
and(p145,a[10],b[4]);
and(p146,a[9],b[5]);
and(p147,a[8],b[6]);
and(p148,a[7],b[7]);
and(p149,a[6],b[8]);
and(p1410,a[5],b[9]);
and(p1411,a[4],b[10]);
and(p1412,a[3],b[11]);
and(p1413,a[2],b[12]);
and(p1414,a[1],b[13]);
and(p1415,a[0],b[14]);
and(p151,a[15],b[0]);
and(p152,a[14],b[1]);
and(p153,a[13],b[2]);
and(p154,a[12],b[3]);
and(p155,a[11],b[4]);
and(p156,a[10],b[5]);
and(p157,a[9],b[6]);
and(p158,a[8],b[7]);
and(p159,a[7],b[8]);
and(p1510,a[6],b[9]);
and(p1511,a[5],b[10]);
and(p1512,a[4],b[11]);
and(p1513,a[3],b[12]);
and(p1514,a[2],b[13]);
and(p1515,a[1],b[14]);
and(p1516,a[0],b[15]);
and(p301,a[15],b[15]);
and(p291,a[15],b[14]);
and(p292,a[14],b[15]);
and(p281,a[15],b[13]);
and(p282,a[14],b[14]);
and(p283,a[13],b[15]);
and(p271,a[15],b[12]);
and(p272,a[14],b[13]);
and(p273,a[13],b[14]);
and(p274,a[12],b[15]);
and(p261,a[15],b[11]);
and(p262,a[14],b[12]);
and(p263,a[13],b[13]);
and(p264,a[12],b[14]);
and(p265,a[11],b[15]);
and(p251,a[15],b[10]);
and(p252,a[14],b[11]);
and(p253,a[13],b[12]);
and(p254,a[12],b[13]);
and(p255,a[11],b[14]);
and(p256,a[10],b[15]);
and(p241,a[15],b[9]);
and(p242,a[14],b[10]);
and(p243,a[13],b[11]);
and(p244,a[12],b[12]);
and(p245,a[11],b[13]);
and(p246,a[10],b[14]);
and(p247,a[9],b[15]);
and(p231,a[15],b[8]);
and(p232,a[14],b[9]);
and(p233,a[13],b[10]);
and(p234,a[12],b[11]);
and(p235,a[11],b[12]);
and(p236,a[10],b[13]);
and(p237,a[9],b[14]);
and(p238,a[8],b[15]);
and(p221,a[15],b[7]);
and(p222,a[14],b[8]);
and(p223,a[13],b[9]);
and(p224,a[12],b[10]);
and(p225,a[11],b[11]);
and(p226,a[10],b[12]);
and(p227,a[9],b[13]);
and(p228,a[8],b[14]);
and(p229,a[7],b[15]);
and(p211,a[15],b[6]);
and(p212,a[14],b[7]);
and(p213,a[13],b[8]);
and(p214,a[12],b[9]);
and(p215,a[11],b[10]);
and(p216,a[10],b[11]);
and(p217,a[9],b[12]);
and(p218,a[8],b[13]);
and(p219,a[7],b[14]);
and(p2110,a[6],b[15]);
and(p201,a[15],b[5]);
and(p202,a[14],b[6]);
and(p203,a[13],b[7]);
and(p204,a[12],b[8]);
and(p205,a[11],b[9]);
and(p206,a[10],b[10]);
and(p207,a[9],b[11]);
and(p208,a[8],b[12]);
and(p209,a[7],b[13]);
and(p2010,a[6],b[14]);
and(p2011,a[5],b[15]);
and(p191,a[15],b[4]);
and(p192,a[14],b[5]);
and(p193,a[13],b[6]);
and(p194,a[12],b[7]);
and(p195,a[11],b[8]);
and(p196,a[10],b[9]);
and(p197,a[9],b[10]);
and(p198,a[8],b[11]);
and(p199,a[7],b[12]);
and(p1910,a[6],b[13]);
and(p1911,a[5],b[14]);
and(p1912,a[4],b[15]);
and(p181,a[15],b[3]);
and(p182,a[14],b[4]);
and(p183,a[13],b[5]);
and(p184,a[12],b[6]);
and(p185,a[11],b[7]);
and(p186,a[10],b[8]);
and(p187,a[9],b[9]);
and(p188,a[8],b[10]);
and(p189,a[7],b[11]);
and(p1810,a[6],b[12]);
and(p1811,a[5],b[13]);
and(p1812,a[4],b[14]);
and(p1813,a[3],b[15]);
and(p171,a[15],b[2]);
and(p172,a[14],b[3]);
and(p173,a[13],b[4]);
and(p174,a[12],b[5]);
and(p175,a[11],b[6]);
and(p176,a[10],b[7]);
and(p177,a[9],b[8]);
and(p178,a[8],b[9]);
and(p179,a[7],b[10]);
and(p1710,a[6],b[11]);
and(p1711,a[5],b[12]);
and(p1712,a[4],b[13]);
and(p1713,a[3],b[14]);
and(p1714,a[2],b[15]);
and(p161,a[15],b[1]);
and(p162,a[14],b[2]);
and(p163,a[13],b[3]);
and(p164,a[12],b[4]);
and(p165,a[11],b[5]);
and(p166,a[10],b[6]);
and(p167,a[9],b[7]);
and(p168,a[8],b[8]);
and(p169,a[7],b[9]);
and(p1610,a[6],b[10]);
and(p1611,a[5],b[11]);
and(p1612,a[4],b[12]);
and(p1613,a[3],b[13]);
and(p1614,a[2],b[14]);
and(p1615,a[1],b[15]);
Butterfly_Mult_HalfAdder  hin1(s1,c1,p1615,p1614);
Butterfly_Mult_HalfAdder  hin2(s2,c2,p1516,p1515);
Butterfly_Mult_FullAdder f1(s1q17,c1q17,c1,p1714,p1713);
Butterfly_Mult_FullAdder f2(s1q16,c1q16,c2,s1,p1613);
Butterfly_Mult_FullAdder f3(s1q15,c1q15,s2,p1514,p1513);
Butterfly_Mult_HalfAdder  h1(s1q14,c1q14,p1415,p1414);
Butterfly_Mult_FullAdder f4(s2q18,c2q18,c1q17,p1813,p1812);
Butterfly_Mult_FullAdder f5(s2q17,c2q17,s1q17,c1q16,p1712);
Butterfly_Mult_FullAdder f6(s2q16,c2q16,s1q16,c1q15,p1612);
Butterfly_Mult_FullAdder f7(s2q15,c2q15,s1q15,c1q14,p1512);
Butterfly_Mult_FullAdder f8(s2q14,c2q14,s1q14,p1413,p1412);
Butterfly_Mult_HalfAdder  h2(s2q13,c2q13,p1314,p1313);
Butterfly_Mult_FullAdder f9(s3q19,c3q19,c2q18,p1912,p1911);
Butterfly_Mult_FullAdder f10(s3q18,c3q18,s2q18,c2q17,p1811);
Butterfly_Mult_FullAdder f11(s3q17,c3q17,s2q17,c2q16,p1711);
Butterfly_Mult_FullAdder f12(s3q16,c3q16,s2q16,c2q15,p1611);
Butterfly_Mult_FullAdder f13(s3q15,c3q15,s2q15,c2q14,p1511);
Butterfly_Mult_FullAdder f14(s3q14,c3q14,s2q14,c2q13,p1411);
Butterfly_Mult_FullAdder f15(s3q13,c3q13,s2q13,p1312,p1311);
Butterfly_Mult_HalfAdder  h3(s3q12,c3q12,p1213,p1212);
Butterfly_Mult_FullAdder f16(s4q20,c4q20,c3q19,p2011,p2010);
Butterfly_Mult_FullAdder f17(s4q19,c4q19,s3q19,c3q18,p1910);
Butterfly_Mult_FullAdder f18(s4q18,c4q18,s3q18,c3q17,p1810);
Butterfly_Mult_FullAdder f19(s4q17,c4q17,s3q17,c3q16,p1710);
Butterfly_Mult_FullAdder f20(s4q16,c4q16,s3q16,c3q15,p1610);
Butterfly_Mult_FullAdder f21(s4q15,c4q15,s3q15,c3q14,p1510);
Butterfly_Mult_FullAdder f22(s4q14,c4q14,s3q14,c3q13,p1410);
Butterfly_Mult_FullAdder f23(s4q13,c4q13,s3q13,c3q12,p1310);
Butterfly_Mult_FullAdder f24(s4q12,c4q12,s3q12,p1211,p1210);
Butterfly_Mult_HalfAdder  h4(s4q11,c4q11,p1112,p1111);
Butterfly_Mult_FullAdder f25(s5q21,c5q21,c4q20,p2110,p219);
Butterfly_Mult_FullAdder f26(s5q20,c5q20,s4q20,c4q19,p209);
Butterfly_Mult_FullAdder f27(s5q19,c5q19,s4q19,c4q18,p199);
Butterfly_Mult_FullAdder f28(s5q18,c5q18,s4q18,c4q17,p189);
Butterfly_Mult_FullAdder f29(s5q17,c5q17,s4q17,c4q16,p179);
Butterfly_Mult_FullAdder f30(s5q16,c5q16,s4q16,c4q15,p169);
Butterfly_Mult_FullAdder f31(s5q15,c5q15,s4q15,c4q14,p159);
Butterfly_Mult_FullAdder f32(s5q14,c5q14,s4q14,c4q13,p149);
Butterfly_Mult_FullAdder f33(s5q13,c5q13,s4q13,c4q12,p139);
Butterfly_Mult_FullAdder f34(s5q12,c5q12,s4q12,c4q11,p129);
Butterfly_Mult_FullAdder f35(s5q11,c5q11,s4q11,p1110,p119);
Butterfly_Mult_HalfAdder  h5(s5q10,c5q10,p1011,p1010);
Butterfly_Mult_FullAdder f36(s6q22,c6q22,c5q21,p229,p228);
Butterfly_Mult_FullAdder f37(s6q21,c6q21,s5q21,c5q20,p218);
Butterfly_Mult_FullAdder f38(s6q20,c6q20,s5q20,c5q19,p208);
Butterfly_Mult_FullAdder f39(s6q19,c6q19,s5q19,c5q18,p198);
Butterfly_Mult_FullAdder f40(s6q18,c6q18,s5q18,c5q17,p188);
Butterfly_Mult_FullAdder f41(s6q17,c6q17,s5q17,c5q16,p178);
Butterfly_Mult_FullAdder f42(s6q16,c6q16,s5q16,c5q15,p168);
Butterfly_Mult_FullAdder f43(s6q15,c6q15,s5q15,c5q14,p158);
Butterfly_Mult_FullAdder f44(s6q14,c6q14,s5q14,c5q13,p148);
Butterfly_Mult_FullAdder f45(s6q13,c6q13,s5q13,c5q12,p138);
Butterfly_Mult_FullAdder f46(s6q12,c6q12,s5q12,c5q11,p128);
Butterfly_Mult_FullAdder f47(s6q11,c6q11,s5q11,c5q10,p118);
Butterfly_Mult_FullAdder f48(s6q10,c6q10,s5q10,p109,p108);
Butterfly_Mult_HalfAdder  h6(s6q9,c6q9,p910,p99);
Butterfly_Mult_FullAdder f49(s7q23,c7q23,c6q22,p238,p237);
Butterfly_Mult_FullAdder f50(s7q22,c7q22,s6q22,c6q21,p227);
Butterfly_Mult_FullAdder f51(s7q21,c7q21,s6q21,c6q20,p217);
Butterfly_Mult_FullAdder f52(s7q20,c7q20,s6q20,c6q19,p207);
Butterfly_Mult_FullAdder f53(s7q19,c7q19,s6q19,c6q18,p197);
Butterfly_Mult_FullAdder f54(s7q18,c7q18,s6q18,c6q17,p187);
Butterfly_Mult_FullAdder f55(s7q17,c7q17,s6q17,c6q16,p177);
Butterfly_Mult_FullAdder f56(s7q16,c7q16,s6q16,c6q15,p167);
Butterfly_Mult_FullAdder f57(s7q15,c7q15,s6q15,c6q14,p157);
Butterfly_Mult_FullAdder f58(s7q14,c7q14,s6q14,c6q13,p147);
Butterfly_Mult_FullAdder f59(s7q13,c7q13,s6q13,c6q12,p137);
Butterfly_Mult_FullAdder f60(s7q12,c7q12,s6q12,c6q11,p127);
Butterfly_Mult_FullAdder f61(s7q11,c7q11,s6q11,c6q10,p117);
Butterfly_Mult_FullAdder f62(s7q10,c7q10,s6q10,c6q9,p107);
Butterfly_Mult_FullAdder f63(s7q9,c7q9,s6q9,p98,p97);
Butterfly_Mult_HalfAdder  h7(s7q8,c7q8,p89,p88);
Butterfly_Mult_FullAdder f64(s8q24,c8q24,c7q23,p247,p246);
Butterfly_Mult_FullAdder f65(s8q23,c8q23,s7q23,c7q22,p236);
Butterfly_Mult_FullAdder f66(s8q22,c8q22,s7q22,c7q21,p226);
Butterfly_Mult_FullAdder f67(s8q21,c8q21,s7q21,c7q20,p216);
Butterfly_Mult_FullAdder f68(s8q20,c8q20,s7q20,c7q19,p206);
Butterfly_Mult_FullAdder f69(s8q19,c8q19,s7q19,c7q18,p196);
Butterfly_Mult_FullAdder f70(s8q18,c8q18,s7q18,c7q17,p186);
Butterfly_Mult_FullAdder f71(s8q17,c8q17,s7q17,c7q16,p176);
Butterfly_Mult_FullAdder f72(s8q16,c8q16,s7q16,c7q15,p166);
Butterfly_Mult_FullAdder f73(s8q15,c8q15,s7q15,c7q14,p156);
Butterfly_Mult_FullAdder f74(s8q14,c8q14,s7q14,c7q13,p146);
Butterfly_Mult_FullAdder f75(s8q13,c8q13,s7q13,c7q12,p136);
Butterfly_Mult_FullAdder f76(s8q12,c8q12,s7q12,c7q11,p126);
Butterfly_Mult_FullAdder f77(s8q11,c8q11,s7q11,c7q10,p116);
Butterfly_Mult_FullAdder f78(s8q10,c8q10,s7q10,c7q9,p106);
Butterfly_Mult_FullAdder f79(s8q9,c8q9,s7q9,c7q8,p96);
Butterfly_Mult_FullAdder f80(s8q8,c8q8,s7q8,p87,p86);
Butterfly_Mult_HalfAdder  h8(s8q7,c8q7,p78,p77);
Butterfly_Mult_FullAdder f81(s9q25,c9q25,c8q24,p256,p255);
Butterfly_Mult_FullAdder f82(s9q24,c9q24,s8q24,c8q23,p245);
Butterfly_Mult_FullAdder f83(s9q23,c9q23,s8q23,c8q22,p235);
Butterfly_Mult_FullAdder f84(s9q22,c9q22,s8q22,c8q21,p225);
Butterfly_Mult_FullAdder f85(s9q21,c9q21,s8q21,c8q20,p215);
Butterfly_Mult_FullAdder f86(s9q20,c9q20,s8q20,c8q19,p205);
Butterfly_Mult_FullAdder f87(s9q19,c9q19,s8q19,c8q18,p195);
Butterfly_Mult_FullAdder f88(s9q18,c9q18,s8q18,c8q17,p185);
Butterfly_Mult_FullAdder f89(s9q17,c9q17,s8q17,c8q16,p175);
Butterfly_Mult_FullAdder f90(s9q16,c9q16,s8q16,c8q15,p165);
Butterfly_Mult_FullAdder f91(s9q15,c9q15,s8q15,c8q14,p155);
Butterfly_Mult_FullAdder f92(s9q14,c9q14,s8q14,c8q13,p145);
Butterfly_Mult_FullAdder f93(s9q13,c9q13,s8q13,c8q12,p135);
Butterfly_Mult_FullAdder f94(s9q12,c9q12,s8q12,c8q11,p125);
Butterfly_Mult_FullAdder f95(s9q11,c9q11,s8q11,c8q10,p115);
Butterfly_Mult_FullAdder f96(s9q10,c9q10,s8q10,c8q9,p105);
Butterfly_Mult_FullAdder f97(s9q9,c9q9,s8q9,c8q8,p95);
Butterfly_Mult_FullAdder f98(s9q8,c9q8,s8q8,c8q7,p85);
Butterfly_Mult_FullAdder f99(s9q7,c9q7,s8q7,p76,p75);
Butterfly_Mult_HalfAdder  h9(s9q6,c9q6,p67,p66);
Butterfly_Mult_FullAdder f100(s10q26,c10q26,c9q25,p265,p264);
Butterfly_Mult_FullAdder f101(s10q25,c10q25,s9q25,c9q24,p254);
Butterfly_Mult_FullAdder f102(s10q24,c10q24,s9q24,c9q23,p244);
Butterfly_Mult_FullAdder f103(s10q23,c10q23,s9q23,c9q22,p234);
Butterfly_Mult_FullAdder f104(s10q22,c10q22,s9q22,c9q21,p224);
Butterfly_Mult_FullAdder f105(s10q21,c10q21,s9q21,c9q20,p214);
Butterfly_Mult_FullAdder f106(s10q20,c10q20,s9q20,c9q19,p204);
Butterfly_Mult_FullAdder f107(s10q19,c10q19,s9q19,c9q18,p194);
Butterfly_Mult_FullAdder f108(s10q18,c10q18,s9q18,c9q17,p184);
Butterfly_Mult_FullAdder f109(s10q17,c10q17,s9q17,c9q16,p174);
Butterfly_Mult_FullAdder f110(s10q16,c10q16,s9q16,c9q15,p164);
Butterfly_Mult_FullAdder f111(s10q15,c10q15,s9q15,c9q14,p154);
Butterfly_Mult_FullAdder f112(s10q14,c10q14,s9q14,c9q13,p144);
Butterfly_Mult_FullAdder f113(s10q13,c10q13,s9q13,c9q12,p134);
Butterfly_Mult_FullAdder f114(s10q12,c10q12,s9q12,c9q11,p124);
Butterfly_Mult_FullAdder f115(s10q11,c10q11,s9q11,c9q10,p114);
Butterfly_Mult_FullAdder f116(s10q10,c10q10,s9q10,c9q9,p104);
Butterfly_Mult_FullAdder f117(s10q9,c10q9,s9q9,c9q8,p94);
Butterfly_Mult_FullAdder f118(s10q8,c10q8,s9q8,c9q7,p84);
Butterfly_Mult_FullAdder f119(s10q7,c10q7,s9q7,c9q6,p74);
Butterfly_Mult_FullAdder f120(s10q6,c10q6,s9q6,p65,p64);
Butterfly_Mult_HalfAdder  h10(s10q5,c10q5,p56,p55);
Butterfly_Mult_FullAdder f121(s11q27,c11q27,c10q26,p274,p273);
Butterfly_Mult_FullAdder f122(s11q26,c11q26,s10q26,c10q25,p263);
Butterfly_Mult_FullAdder f123(s11q25,c11q25,s10q25,c10q24,p253);
Butterfly_Mult_FullAdder f124(s11q24,c11q24,s10q24,c10q23,p243);
Butterfly_Mult_FullAdder f125(s11q23,c11q23,s10q23,c10q22,p233);
Butterfly_Mult_FullAdder f126(s11q22,c11q22,s10q22,c10q21,p223);
Butterfly_Mult_FullAdder f127(s11q21,c11q21,s10q21,c10q20,p213);
Butterfly_Mult_FullAdder f128(s11q20,c11q20,s10q20,c10q19,p203);
Butterfly_Mult_FullAdder f129(s11q19,c11q19,s10q19,c10q18,p193);
Butterfly_Mult_FullAdder f130(s11q18,c11q18,s10q18,c10q17,p183);
Butterfly_Mult_FullAdder f131(s11q17,c11q17,s10q17,c10q16,p173);
Butterfly_Mult_FullAdder f132(s11q16,c11q16,s10q16,c10q15,p163);
Butterfly_Mult_FullAdder f133(s11q15,c11q15,s10q15,c10q14,p153);
Butterfly_Mult_FullAdder f134(s11q14,c11q14,s10q14,c10q13,p143);
Butterfly_Mult_FullAdder f135(s11q13,c11q13,s10q13,c10q12,p133);
Butterfly_Mult_FullAdder f136(s11q12,c11q12,s10q12,c10q11,p123);
Butterfly_Mult_FullAdder f137(s11q11,c11q11,s10q11,c10q10,p113);
Butterfly_Mult_FullAdder f138(s11q10,c11q10,s10q10,c10q9,p103);
Butterfly_Mult_FullAdder f139(s11q9,c11q9,s10q9,c10q8,p93);
Butterfly_Mult_FullAdder f140(s11q8,c11q8,s10q8,c10q7,p83);
Butterfly_Mult_FullAdder f141(s11q7,c11q7,s10q7,c10q6,p73);
Butterfly_Mult_FullAdder f142(s11q6,c11q6,s10q6,c10q5,p63);
Butterfly_Mult_FullAdder f143(s11q5,c11q5,s10q5,p54,p53);
Butterfly_Mult_HalfAdder  h11(s11q4,c11q4,p45,p44);
Butterfly_Mult_FullAdder f144(s12q28,c12q28,c11q27,p283,p282);
Butterfly_Mult_FullAdder f145(s12q27,c12q27,s11q27,c11q26,p272);
Butterfly_Mult_FullAdder f146(s12q26,c12q26,s11q26,c11q25,p262);
Butterfly_Mult_FullAdder f147(s12q25,c12q25,s11q25,c11q24,p252);
Butterfly_Mult_FullAdder f148(s12q24,c12q24,s11q24,c11q23,p242);
Butterfly_Mult_FullAdder f149(s12q23,c12q23,s11q23,c11q22,p232);
Butterfly_Mult_FullAdder f150(s12q22,c12q22,s11q22,c11q21,p222);
Butterfly_Mult_FullAdder f151(s12q21,c12q21,s11q21,c11q20,p212);
Butterfly_Mult_FullAdder f152(s12q20,c12q20,s11q20,c11q19,p202);
Butterfly_Mult_FullAdder f153(s12q19,c12q19,s11q19,c11q18,p192);
Butterfly_Mult_FullAdder f154(s12q18,c12q18,s11q18,c11q17,p182);
Butterfly_Mult_FullAdder f155(s12q17,c12q17,s11q17,c11q16,p172);
Butterfly_Mult_FullAdder f156(s12q16,c12q16,s11q16,c11q15,p162);
Butterfly_Mult_FullAdder f157(s12q15,c12q15,s11q15,c11q14,p152);
Butterfly_Mult_FullAdder f158(s12q14,c12q14,s11q14,c11q13,p142);
Butterfly_Mult_FullAdder f159(s12q13,c12q13,s11q13,c11q12,p132);
Butterfly_Mult_FullAdder f160(s12q12,c12q12,s11q12,c11q11,p122);
Butterfly_Mult_FullAdder f161(s12q11,c12q11,s11q11,c11q10,p112);
Butterfly_Mult_FullAdder f162(s12q10,c12q10,s11q10,c11q9,p102);
Butterfly_Mult_FullAdder f163(s12q9,c12q9,s11q9,c11q8,p92);
Butterfly_Mult_FullAdder f164(s12q8,c12q8,s11q8,c11q7,p82);
Butterfly_Mult_FullAdder f165(s12q7,c12q7,s11q7,c11q6,p72);
Butterfly_Mult_FullAdder f166(s12q6,c12q6,s11q6,c11q5,p62);
Butterfly_Mult_FullAdder f167(s12q5,c12q5,s11q5,c11q4,p52);
Butterfly_Mult_FullAdder f168(s12q4,c12q4,s11q4,p43,p42);
Butterfly_Mult_HalfAdder  h12(s12q3,c12q3,p34,p33);
Butterfly_Mult_FullAdder f169(s13q29,c13q29,c12q28,p292,p291);
Butterfly_Mult_FullAdder f170(s13q28,c13q28,s12q28,c12q27,p281);
Butterfly_Mult_FullAdder f171(s13q27,c13q27,s12q27,c12q26,p271);
Butterfly_Mult_FullAdder f172(s13q26,c13q26,s12q26,c12q25,p261);
Butterfly_Mult_FullAdder f173(s13q25,c13q25,s12q25,c12q24,p251);
Butterfly_Mult_FullAdder f174(s13q24,c13q24,s12q24,c12q23,p241);
Butterfly_Mult_FullAdder f175(s13q23,c13q23,s12q23,c12q22,p231);
Butterfly_Mult_FullAdder f176(s13q22,c13q22,s12q22,c12q21,p221);
Butterfly_Mult_FullAdder f177(s13q21,c13q21,s12q21,c12q20,p211);
Butterfly_Mult_FullAdder f178(s13q20,c13q20,s12q20,c12q19,p201);
Butterfly_Mult_FullAdder f179(s13q19,c13q19,s12q19,c12q18,p191);
Butterfly_Mult_FullAdder f180(s13q18,c13q18,s12q18,c12q17,p181);
Butterfly_Mult_FullAdder f181(s13q17,c13q17,s12q17,c12q16,p171);
Butterfly_Mult_FullAdder f182(s13q16,c13q16,s12q16,c12q15,p161);
Butterfly_Mult_FullAdder f183(s13q15,c13q15,s12q15,c12q14,p151);
Butterfly_Mult_FullAdder f184(s13q14,c13q14,s12q14,c12q13,p141);
Butterfly_Mult_FullAdder f185(s13q13,c13q13,s12q13,c12q12,p131);
Butterfly_Mult_FullAdder f186(s13q12,c13q12,s12q12,c12q11,p121);
Butterfly_Mult_FullAdder f187(s13q11,c13q11,s12q11,c12q10,p111);
Butterfly_Mult_FullAdder f188(s13q10,c13q10,s12q10,c12q9,p101);
Butterfly_Mult_FullAdder f189(s13q9,c13q9,s12q9,c12q8,p91);
Butterfly_Mult_FullAdder f190(s13q8,c13q8,s12q8,c12q7,p81);
Butterfly_Mult_FullAdder f191(s13q7,c13q7,s12q7,c12q6,p71);
Butterfly_Mult_FullAdder f192(s13q6,c13q6,s12q6,c12q5,p61);
Butterfly_Mult_FullAdder f193(s13q5,c13q5,s12q5,c12q4,p51);
Butterfly_Mult_FullAdder f194(s13q4,c13q4,s12q4,c12q3,p41);
Butterfly_Mult_FullAdder f195(s13q3,c13q3,s12q3,p32,p31);
Butterfly_Mult_HalfAdder  h13(s13q2,c13q2,p23,p22);
assign x={p301,s13q29,s13q28,s13q27,s13q26,s13q25,s13q24,s13q23,s13q22,s13q21,s13q20,s13q19,s13q18,s13q17,s13q16,s13q15,s13q14,s13q13,s13q12,s13q11,s13q10,s13q9,s13q8,s13q7,s13q6,s13q5,s13q4,s13q3,p21,p11};
assign y={c13q29,c13q28,c13q27,c13q26,c13q25,c13q24,c13q23,c13q22,c13q21,c13q20,c13q19,c13q18,c13q17,c13q16,c13q15,c13q14,c13q13,c13q12,c13q11,c13q10,c13q9,c13q8,c13q7,c13q6,c13q5,c13q4,c13q3,c13q2,s13q2,p12};
Butterfly_Mult_Wallace_Adder wadd001(z,t,x,y);
assign prod={t,z,p01};
endmodule
